//INV for use in these modules
module not1 (in1,out);
input in1;
output out;
assign out = ~in1;
endmodule


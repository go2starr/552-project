/* se11_16.v - 11 to 16-bit sign extender */
module se8_16(
	      // Inputs
	      in,
	      // Outputs
	      out
	      );
   // Inputs
   input [10:0] in;

   // Outputs
   output [15:0] out;
endmodule // se8_16



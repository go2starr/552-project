/* se8_16.v - 8 to 16-bit sign extender */
module se8_16(
	      // Inputs
	      in,
	      // Outputs
	      out
	      );
   // Inputs
   input [7:0] in;

   // Outputs
   output [15:0] out;
endmodule // se8_16


`include "testbench.v"

`define DEBUG 1

// t_proc_bench.v
module t_proc_bench();
   // DUT Outputs
   wire err;

   // Clkrst
   wire clk, rst;
   clkrst cr(clk, rst, err);
   
   // CPU - DUT
   proc dut (.clk(clk),
             .rst(rst),
             .err(err)
             );


   // Counters
   integer i,j,k, no_errs;


   initial begin
      `info("Starting tests");

      /****************************************
       *  Check reset conditions
       *****************************************/
      `tic;
      `test(0, dut.pc, "PC did not reset to 0");


      `tic;
      `tic;


      /****************************************
       *  Test first instruction
       ****************************************/
      `info("lbi r0, 0x10");

      $display("PC: %h \t Instr: %h", dut.pc, dut.instr);
      // dut
      `test(16'h c010, dut.instr, "Instruction does not match: lbi r0, 0x10");
      `test(16'h 0, dut.pc, "PC should be 0 on start");
      `test(16'h 10, dut.alu.Out, "ALU output should be zero");

      // aopd
      `test(16'h 10, dut.aopd.opB, "ALU op decode output should be 0x10");
      `test(16'h c010, dut.aopd.instr, "Input to alu_op_decode should be instruction");
      `test(7'b 1100000, dut.aopd.op, "Op should be correct");

      // alu
      `test(16'h 10, dut.alu.opB, "ALU opB should be 0x10");
      `test(16'h 10, dut.alu.B, "ALU input should be 0x10 (immediate value)");
      `test(5'd  19, dut.alu.Op, "ALU op should be LBI");
      `test(16'h 10, dut.alu.Out, "ALU output should be 0x10");

      // add (destination decode)
      `test(16'h c010, dut.add.instr, "add instruction should be correct");
      `test(3'h  0,    dut.add.rd, "add register select should be zero");
      
      // write to rf
      `test(16'h 0, dut.rf_ws, "RF write select should be zero");
      `test(16'h 10, dut.rf_wd, "RF write data should be 0x10");
      
      /****************************************/
      `tic;
      /****************************************/
      `test(16'h10, dut.rf.rf0.my_regs0.q, "R0 does not contain 0x10 after a lbi 0x10");

      // dut
      `test(16'h c101, dut.instr, "Instruction does not match: lbi r1, 0x01");
      `test(16'h 2, dut.pc, "PC should be 2 after first instruction");

      // add (destination decode)
      
      // write to rf
      `test(16'h 01, dut.rf_ws, "RF write select should be one");      
      `test(16'h 01, dut.rf_wd, "RF write data should be 0x01");

      

      /****************************************/
      `tic;
      /****************************************/
      `test(16'h01, dut.rf.rf0.my_regs1.q, "R1 does not contain 0x01 after lbi r1, 0x01");

      `info("add r2, r0, r1");

      // dut
      `test(16'h 4, dut.pc, "PC should be 4 after second instruction");
      `test(16'h d828, dut.instr, "Instruction does not match: add r2, r0, r1");

      // rf
      `test(3'h 0, dut.rf.read1regsel, "RF internal read1 select is not 0");
      `test(3'h 1, dut.rf.read2regsel, "RF internal read2 select is not 1");      
      `test(16'h 10, dut.rf.read1data, "RF read1 data is not 0x10");
      `test(16'h 01, dut.rf.read2data, "RF read2 data is not 0x10");      
      
      `test(16'h 10, dut.rf.rf0.my_regs0.q, "RF did not hold value(0x10) for r0");
      `test(16'h 01, dut.rf.rf0.my_regs1.q, "RF did not hold value(0x01) for r1");      
      
      
      `test(3'h 0, dut.rf_rs1, "RF select 1 is not r0");
      `test(3'h 1, dut.rf_rs2, "RF select 2 is not r1");
      `test(3'h 10, dut.rf_rd1, "RF data 1 is not 0x10");
      `test(3'h 1, dut.rf_rd2, "RF data 2 is not 0x1");      
      
      

      // alu
      `test(16'h 10, dut.alu.A, "ALU primary op is not 0x10");
      `test(16'h 01, dut.alu.B, "ALU primary op is not 0x01");      
      
      `test(16'h 11, dut.alu.Out, "ALU output is not 0x11");

      // result
      `test(16'h 11, dut.rf.rf0.my_regs2.q, "R0(0x10) + R1(0x01) not put into R2");

      

      `info("Tests complete");
      $finish;
   end   

endmodule // t_proc_bench


/* se5_16.v - 5 to 16-bit sign extender */
module se5_16(
	      // Inputs
	      in,
	      // Outputs
	      out
	      );
   // Inputs
   input [4:0] in;

   // Outputs
   output [15:0] out;
endmodule // se5_16
